//////////////////////////////////////////////////////////////////////////////////
//
// VGA Driver Controller
//
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps
`include "Display640x480.vh"

module pong(
    input clock,
    output reg [3:0] red,
    output reg [3:0] green,
    output reg [3:0] blue,
    output hsync, vsync, avideo,
    input switch,
    input reset,
    input pushUp,
    input pushDown
  );

   wire [`xbits-1:0] x;
   wire [`ybits-1:0] y;
   wire [9:0] y_I_Barra;
   wire [9:0] y_S_Barra;
   wire [9:0] x_I_Bola;
   wire [9:0] x_F_Bola;
   wire [9:0] y_S_Bola;
   wire [9:0] y_I_Bola;
   wire activevideo;
   wire sentido;

   reg aux_reset = 0;
   reg aux_reset1 = 0;

  assign avideo = activevideo;

  reg [1:0] clock_count = 0;
  always @(posedge clock) begin : proc_clock_count
    clock_count <= clock_count + 2'b01;
  end

  MOVBarra myMov
  (
    clock, 
    reset, 
    pushUp, 
    pushDown, 
    y_S_Barra, 
    y_I_Barra,
    aux_reset
  );
   
  impact impact
  (
    .clock(clock),
    .reset(reset),
    .Pos_barra_y_S(y_S_Barra),
    .Pos_barra_y_I(y_I_Barra),
    .Pos_bola_I_x(x_I_Bola),
    .Pos_bola_F_x(x_F_Bola),
    .Pos_bola_S_y(y_S_Bola),
    .Pos_bola_I_y(y_I_Bola),
    .sentido_x(sentido),
    .ponto(ponto),
    .setor1(setor1),
    .setor2(setor2),
    .setor3(setor3),
    .setor4(setor4),
    .setor5(setor5),
    .setor6(setor6)
  );

  MOVBola myMovBola
  (
    clock, 
    reset,
    sentido,
    x_F_Bola, 
    x_I_Bola,
    y_S_Bola,
    y_I_Bola,
    Pos_barra_y_S,
    Pos_barra_y_I,
    ponto, 
    setor1,
    setor2,
    setor3,
    setor4,
    setor5,
    setor6,
    aux_reset
  );

  VGASyncTimer myVGATimer
  (
    clock, 
    hsync, 
    vsync, 
    activevideo, 
    x, 
    y
  );

  always @(posedge clock) begin
    //desenho menu
    if (switch == 0) begin

      aux_reset <= 0;
      aux_reset1 <= 0;

      red[3:0] <= (activevideo == 1) ? (  
                                        ((x>=200 && x<=204) && (y>=80 && y<=135)) || ((y>=80 && y<=84) && (x>=204 && x<=232)) || ((y>=80 && y<=109) && (x>=232 && x<=236)) || ((y>=105 && y<=109) && (x>=204 && x<=232)) ||
                                        ((x>=256 && x<=260) && (y>=80 && y<=135)) || ((y>=80 && y<=84) && (x>=260 && x<=288)) || ((y>=80 && y<=135) && (x>=288 && x<=292)) || ((y>=131 && y<=135) && (x>=260 && x<=288)) ||
                                        ((x>=308 && x<=312) && (y>=80 && y<=135)) || ((y>=80 && y<=135) && (x>=340 && x<=344))|| ((y>=80 && y<=84) && (x>=312 && x<=316)) || ((y>=84 && y<=88) && (x>=316 && x<=320))  || ((y>=88 && y<=92) && (x>=320 && x<=324)) || ((y>=92 && y<=96) && (x>=324 && x<=328)) || ((y>=96 && y<=100) && (x>=328 && x<=332)) || ((y>=100 && y<=104) && (x>=332 && x<=336)) || ((y>=104 && y<=108) && (x>=336 && x<=340)) ||
                                        ((x>=364 && x<=368) && (y>=80 && y<=135)) || ((y>=80 && y<=84) && (x>=368 && x<=394)) || ((y>=106 && y<=135) && (x>=392 && x<=396)) || ((y>=131 && y<=135) && (x>=368 && x<=394)) || ((y>=106 && y<=110) && (x>=380 && x<=394)) ||
                                        ((x>=30 && x<=33) && (y>=210 && y<=250)) || ((x>=100 && x<=104) && (y>=210 && y<=216)) || ((x>=200 && x<=204) && (y>=310 && y<=316)) || ((x>=300 && x<=304) && (y>=250 && y<=256)) ||
                                        ((x>=318 && x<=322) && (y>=420 && y<=450)) || ((y>=446 && y<=450) && (x>=322 && x<=342)) || ((x>=342 && x<=346) && (y>=420 && y<=450)) || ((y>=430 && y<=433) && (x>=327 && x<=337)) || ((x>=331 && x<=333) && (y>=410 && y<=433)) || ((x>=310 && x<=311) && (y>=410 && y<=423)) || ((x>=307 && x<=311) && (y>=444 && y<=450))
      ? 4'b1111 : 4'b0000) : (4'b0);
      
      blue[3:0] <= (activevideo == 1) ? (((x>=394 && x<=398) && (y>=150 && y<=180)) || ((y>=150 && y<=154) && (x>=398 && x<=413)) || ((y>=160 && y<=164) && (x>=398 && x<=413)) ||
                                        ((x>=423 && x<=427) && (y>=150 && y<=180)) || ((y>=150 && y<=154) && (x>=427 && x<=442)) ||  ((x>=438 && x<=442) && (y>=150 && y<=164)) || ((y>=165 && y<=169) && (x>=427 && x<=442)) ||                                               
                                        ((x>=452 && x<=456) && (y>=150 && y<=180)) || ((y>=150 && y<=154) && (x>=456 && x<=471)) ||  ((x>=467 && x<=471) && (y>=170 && y<=180)) || ((y>=166 && y<=170) && (x>=465 && x<=471)) || ((y>=176 && y<=180) && (x>=456 && x<=471)) ||
                                        ((x>=481 && x<=485) && (y>=150 && y<=180)) || ((y>=150 && y<=154) && (x>=485 && x<=500)) ||  ((x>=496 && x<=500) && (y>=150 && y<=180)) || ((y>=165 && y<=169) && (x>=485 && x<=500)) ||
                                        ((x>=30 && x<=33) && (y>=210 && y<=250)) || ((x>=100 && x<=104) && (y>=210 && y<=216)) || ((x>=200 && x<=204) && (y>=310 && y<=316)) || ((x>=300 && x<=304) && (y>=250 && y<=256)) ||
                                        ((x>=318 && x<=322) && (y>=420 && y<=450)) || ((y>=446 && y<=450) && (x>=322 && x<=342)) || ((x>=342 && x<=346) && (y>=420 && y<=450)) || ((y>=430 && y<=433) && (x>=327 && x<=337)) || ((x>=331 && x<=333) && (y>=410 && y<=433)) || ((x>=310 && x<=311) && (y>=410 && y<=423)) || ((x>=307 && x<=311) && (y>=444 && y<=450))
       ? 4'b1111 : 4'b0000) : (4'b0);
      
      green[3:0] <= (activevideo == 1) ?  (
                                          ((x>=30 && x<=33) && (y>=210 && y<=250)) || ((x>=100 && x<=104) && (y>=210 && y<=216)) || ((x>=200 && x<=204) && (y>=310 && y<=316)) || ((x>=300 && x<=304) && (y>=250 && y<=256)) ||
                                          ((x>=318 && x<=322) && (y>=420 && y<=450)) || ((y>=446 && y<=450) && (x>=322 && x<=342)) || ((x>=342 && x<=346) && (y>=420 && y<=450)) || ((y>=430 && y<=433) && (x>=327 && x<=337)) || ((x>=331 && x<=333) && (y>=410 && y<=433)) || ((x>=310 && x<=311) && (y>=410 && y<=423)) || ((x>=307 && x<=311) && (y>=444 && y<=450))
     ? 4'b1111 : 4'b0000) : (4'b0);
      
    end
  
    else begin
      
      if (aux_reset == 0 && aux_reset1 == 0)
        aux_reset <= 1;

      if(aux_reset == 1 && aux_reset1 == 0) begin
        aux_reset1 <= 1;
        aux_reset <= 0;
      end

      red[3:0] <= (activevideo == 1) ?  (
                                        ((y>=4 && y<=20) && (x>=15 && x<=16)) || ((y>=4 && y<=5) && (x>=17 && x<=21)) || ((y>=4 && y<=8) && (x>=21 && x<=22)) || ((y>=9 && y<=10) && (x>=17 && x<=22)) ||
                                        ((x>=318 && x<=322) && (y>=0 && y<=25)) ||
                                        ((y>=25 && y<=28) || y>=476 || (x>=636 && y>=25)) || ((x>=30 && x<=33) && (y>=y_S_Barra && y<=y_I_Barra)) || ( (x>=x_I_Bola && x<=x_F_Bola) && (y>=y_S_Bola && y<=y_I_Bola)) ? 4'b1111 : 4'b0000) : (4'b0);

      blue[3:0] <= (activevideo == 1) ? (
                                        ((x>=318 && x<=322) && (y>=0 && y<=25)) ||
                                        ((y>=25 && y<=28) || y>=476 || (x>=636 && y>=25)) || ((x>=30 && x<=33) && (y>=y_S_Barra && y<=y_I_Barra)) || ((x>=x_I_Bola && x<=x_F_Bola) && (y>=y_S_Bola && y<=y_I_Bola)) ? 4'b1111 : 4'b0000) : (4'b0);
      
      green[3:0] <= (activevideo == 1) ?  (
                                          ((x>=318 && x<=322) && (y>=0 && y<=25)) ||
                                          ((y>=4 && y<=20) && (x>=336 && x<=337)) || ((y>=4 && y<=5) && (x>=337 && x<=347)) || ((y>=19 && y<=20) && (x>=337 && x<=347)) ||
                                          ((y>=25 && y<=28) || y>=476 || (x>=636 && y>=25)) || ((x>=30 && x<=33) && (y>=y_S_Barra && y<=y_I_Barra)) || ((x>=x_I_Bola && x<=x_F_Bola) && (y>=y_S_Bola && y<=y_I_Bola)) ? 4'b1111 : 4'b0000) : (4'b0);
    end
  end

endmodule